module multiply(a, b, c, cout, acc); 
	input[7:0] a; 
	input[7:0] b; 
	input[7:0] acc; 
	output[15:0] cout; 
	output[15:0] c; 
	assign cout = a*b; 
	assign c = acc +cout; 
endmodule
